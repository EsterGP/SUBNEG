module mem #(
    parameters
) (
    ports
);
    
endmodule