module mem_data #(
    parameters
) (
    ports
);
    
endmodule