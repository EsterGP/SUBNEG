module mem_rom #(
    parameters
) (
    ports
);
    
endmodule